library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity DDS is
    port (
        clk       : in  std_logic;
        reset     : in  std_logic;
        freq_ctrl : in  std_logic_vector(31 downto 0);
        sine_out  : out std_logic_vector(11 downto 0)
    );
end entity DDS;

architecture Behavioral of DDS is

    signal phase_acc      : unsigned(31 downto 0) := (others => '0');
    signal sine_lut_index : unsigned(7 downto 0);

   
    type sine_lut_type is array (0 to 255) of std_logic_vector(11 downto 0);
    
    constant sine_lut : sine_lut_type := 
    (
    "011111111111",
    "100000110001",
    "100001100011",
    "100010010110",
    "100011001000",
    "100011111010",
    "100100101011",
    "100101011101",
    "100110001110",
    "100111000000",
    "100111110000",
    "101000100001",
    "101001010001",
    "101010000001",
    "101010110001",
    "101011100000",
    "101100001110",
    "101100111101",
    "101101101010",
    "101110010111",
    "101111000100",
    "101111110000",
    "110000011011",
    "110001000110",
    "110001110000",
    "110010011010",
    "110011000010",
    "110011101010",
    "110100010010",
    "110100111000",
    "110101011110",
    "110110000010",
    "110110100110",
    "110111001010",
    "110111101100",
    "111000001101",
    "111000101101",
    "111001001101",
    "111001101011",
    "111010001001",
    "111010100101",
    "111011000000",
    "111011011011",
    "111011110100",
    "111100001100",
    "111100100011",
    "111100111001",
    "111101001110",
    "111101100010",
    "111101110101",
    "111110000110",
    "111110010111",
    "111110100110",
    "111110110100",
    "111111000001",
    "111111001100",
    "111111010111",
    "111111100000",
    "111111101000",
    "111111101111",
    "111111110100",
    "111111111000",
    "111111111100",
    "111111111101",
    "111111111110",
    "111111111101",
    "111111111100",
    "111111111000",
    "111111110100",
    "111111101111",
    "111111101000",
    "111111100000",
    "111111010111",
    "111111001100",
    "111111000001",
    "111110110100",
    "111110100110",
    "111110010111",
    "111110000110",
    "111101110101",
    "111101100010",
    "111101001110",
    "111100111001",
    "111100100011",
    "111100001100",
    "111011110100",
    "111011011011",
    "111011000000",
    "111010100101",
    "111010001001",
    "111001101011",
    "111001001101",
    "111000101101",
    "111000001101",
    "110111101100",
    "110111001010",
    "110110100110",
    "110110000010",
    "110101011110",
    "110100111000",
    "110100010010",
    "110011101010",
    "110011000010",
    "110010011010",
    "110001110000",
    "110001000110",
    "110000011011",
    "101111110000",
    "101111000100",
    "101110010111",
    "101101101010",
    "101100111101",
    "101100001110",
    "101011100000",
    "101010110001",
    "101010000001",
    "101001010001",
    "101000100001",
    "100111110000",
    "100111000000",
    "100110001110",
    "100101011101",
    "100100101011",
    "100011111010",
    "100011001000",
    "100010010110",
    "100001100011",
    "100000110001",
    "011111111111",
    "011111001101",
    "011110011011",
    "011101101000",
    "011100110110",
    "011100000100",
    "011011010011",
    "011010100001",
    "011001110000",
    "011000111110",
    "011000001110",
    "010111011101",
    "010110101101",
    "010101111101",
    "010101001101",
    "010100011110",
    "010011110000",
    "010011000001",
    "010010010100",
    "010001100111",
    "010000111010",
    "010000001110",
    "001111100011",
    "001110111000",
    "001110001110",
    "001101100100",
    "001100111100",
    "001100010100",
    "001011101100",
    "001011000110",
    "001010100000",
    "001001111100",
    "001001011000",
    "001000110100",
    "001000010010",
    "000111110001",
    "000111010001",
    "000110110001",
    "000110010011",
    "000101110101",
    "000101011001",
    "000100111110",
    "000100100011",
    "000100001010",
    "000011110010",
    "000011011011",
    "000011000101",
    "000010110000",
    "000010011100",
    "000010001001",
    "000001111000",
    "000001100111",
    "000001011000",
    "000001001010",
    "000000111101",
    "000000110010",
    "000000100111",
    "000000011110",
    "000000010110",
    "000000001111",
    "000000001010",
    "000000000110",
    "000000000010",
    "000000000001",
    "000000000000",
    "000000000001",
    "000000000010",
    "000000000110",
    "000000001010",
    "000000001111",
    "000000010110",
    "000000011110",
    "000000100111",
    "000000110010",
    "000000111101",
    "000001001010",
    "000001011000",
    "000001100111",
    "000001111000",
    "000010001001",
    "000010011100",
    "000010110000",
    "000011000101",
    "000011011011",
    "000011110010",
    "000100001010",
    "000100100011",
    "000100111110",
    "000101011001",
    "000101110101",
    "000110010011",
    "000110110001",
    "000111010001",
    "000111110001",
    "001000010010",
    "001000110100",
    "001001011000",
    "001001111100",
    "001010100000",
    "001011000110",
    "001011101100",
    "001100010100",
    "001100111100",
    "001101100100",
    "001110001110",
    "001110111000",
    "001111100011",
    "010000001110",
    "010000111010",
    "010001100111",
    "010010010100",
    "010011000001",
    "010011110000",
    "010100011110",
    "010101001101",
    "010101111101",
    "010110101101",
    "010111011101",
    "011000001110",
    "011000111110",
    "011001110000",
    "011010100001",
    "011011010011",
    "011100000100",
    "011100110110",
    "011101101000",
    "011110011011",
    "011111001101"
    );
begin
    process (clk, reset)
    begin
        if reset = '0' then
            phase_acc <= (others => '0');
            
        elsif rising_edge(clk) then
            phase_acc <= phase_acc + unsigned(freq_ctrl);
            
            
  
        end if;
    end process;
    sine_lut_index <= phase_acc(31 downto 24); 
    sine_out <= sine_lut(to_integer(sine_lut_index));
   
end architecture Behavioral;
